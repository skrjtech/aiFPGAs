// STSource.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module STSource (
		input  wire        clk,       //       clk.clk
		input  wire        reset,     // clk_reset.reset
		output wire [31:0] src_data,  //       src.data
		output wire [0:0]  src_valid, //          .valid
		input  wire        src_ready  //          .ready
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (0),
		.USE_CHANNEL      (0),
		.USE_ERROR        (0),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (0),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (1),
		.ST_ERROR_W       (1),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (1),
		.VHDL_ID          (0)
	) st_source_bfm_0 (
		.clk               (clk),       //       clk.clk
		.reset             (reset),     // clk_reset.reset
		.src_data          (src_data),  //       src.data
		.src_valid         (src_valid), //          .valid
		.src_ready         (src_ready), //          .ready
		.src_startofpacket (),          // (terminated)
		.src_endofpacket   (),          // (terminated)
		.src_empty         (),          // (terminated)
		.src_channel       (),          // (terminated)
		.src_error         ()           // (terminated)
	);

endmodule
