
module Top #(
    parameter
        
) (
    ports
);
    
endmodule