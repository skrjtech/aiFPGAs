
// Random 
// ------------------------------------------------------------------------------------------------
module Random #(
    parameter
        DWIDTH = 32
) (
    input  wire [DWIDTH - 1: 0] SEED,
    output wire [DWIDTH - 1: 0] OUT
);
/*
Description

    ・　乱数

    Parameter 
        None

    in : SEED   シード値
    out: OUT    出力値
*/

// ?????
// ----------------------------------------------

endmodule