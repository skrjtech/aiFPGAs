// int 4byte to 8byte
// ------------------------------------------------------------------------------------------------
module Int2Long (
    input  wire IN,
    output wire OUT
);
/*
Description

    ・　整数値サイズ大に変換

    Parameter 
        None

    in : IN     入力値
    out: OUT    出力値
*/

// 型変換処理
// ----------------------------------------------
    
endmodule

// Long 8byte to 4byte
// ------------------------------------------------------------------------------------------------
module Long2Int (
    input  wire IN,
    output wire OUT
);
/*
Description

    ・　整数値サイズ小に変換

    Parameter 
        None

    in : IN     入力値
    out: OUT    出力値
*/

// 型変換処理
// ----------------------------------------------

endmodule

// int 4byte to float 4byte
// ------------------------------------------------------------------------------------------------
module Int2Float (
    input  wire IN,
    output wire OUT
);
/*
Description

    ・　整数値から浮動小数点に変換

    Parameter 
        None

    in : IN     入力値
    out: OUT    出力値
*/

// 型変換処理
// ----------------------------------------------

endmodule

// int 4byte to float 8byte
// ------------------------------------------------------------------------------------------------
module Int2FloatLong (
    input  wire IN,
    output wire OUT
);
/*
Description

    ・　整数値から浮動小数点大に変換

    Parameter 
        None

    in : IN     入力値
    out: OUT    出力値
*/

// 型変換処理
// ----------------------------------------------

endmodule

// int 4byte to half float 2byte
// ------------------------------------------------------------------------------------------------
module Int2HalfFloat (
    input  wire IN,
    output wire OUT
);
/*
Description

    ・　整数値から浮動小数点小に変換

    Parameter 
        None

    in : IN     入力値
    out: OUT    出力値
*/

// 型変換処理
// ----------------------------------------------

endmodule

// float 4byte to int 4byte
// ------------------------------------------------------------------------------------------------
module Float2Int (
    input  wire IN,
    output wire OUT
);
/*
Description

    ・　浮動小数点から整数値に変換

    Parameter 
        None

    in : IN     入力値
    out: OUT    出力値
*/

// 型変換処理
// ----------------------------------------------

endmodule

// float 8byte to int 4byte
// ------------------------------------------------------------------------------------------------
module FloatLong2Int (
    input  wire IN,
    output wire OUT
);
/*
Description

    ・　浮動小数点大から整数値に変換

    Parameter 
        None

    in : IN     入力値
    out: OUT    出力値
*/

// 型変換処理
// ----------------------------------------------
    
endmodule

// half float 2byte to int 4byte
// ------------------------------------------------------------------------------------------------
module HalfFloat2Int (
    input  wire IN,
    output wire OUT
);
/*
Description

    ・　浮動小数点小から整数値に変換

    Parameter 
        None

    in : IN     入力値
    out: OUT    出力値
*/

// 型変換処理
// ----------------------------------------------
    
endmodule